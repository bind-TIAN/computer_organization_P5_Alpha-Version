`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:43:54 09/05/2020 
// Design Name: 
// Module Name:    yumen_bgtz 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module yumen_bgtz(
    input a,
    input b,
    output c
    );
	 assign c = a & b;

endmodule
